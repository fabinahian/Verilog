module half_Adder (
    a,
    b,
    carry,
    sum
);

  input a, b;
  output carry, sum;

  


endmodule
