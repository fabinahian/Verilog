module testbench;

initial begin
    $display ("Hello, world!");
end

endmodule